module rho_pi_chi_iota(out, rc, in0, in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, in11, in12, in13, in14, in15, in16, in17, in18, in19, in20, in21, in22, in23, in24);
    input [63:0 ] in0, in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, in11, in12, in13, in14, in15, in16, in17, in18, in19, in20, in21, in22, in23, in24;
    input [7:0]   rc;
    output [1599:0] out;
    
    wire [63:0] reg0_iota, reg0_chi;

    assign reg0_chi = ~({in6 [43:0],in6 [63:44]}) & {in12[42:0],in12[63:43]};

    assign  {reg0_iota[0], reg0_iota[32], reg0_iota[48], reg0_iota[56], reg0_iota[60], reg0_iota[61], reg0_iota[62], reg0_iota[63]} = 
            {in0[0],       in0[32],       in0[48],       in0[56],       in0[60],       in0[61],       in0[62],       in0[63]} ^ rc[7:0];

    assign  {reg0_iota[59:57] , reg0_iota[55:49], reg0_iota[47:33], reg0_iota[31:1]} = 
            {in0[59:57],        in0[55:49],       in0[47:33],       in0[31:1]};

    // assign out[1599:1536] = in0                      ^ (~({in6 [43:0],in6 [63:44]}) & {in12[42:0],in12[63:43]});
    assign out[1599:1536] = reg0_iota                ^ reg0_chi;
    assign out[1535:1472] = {in6 [43:0],in6 [63:44]} ^ (~({in12[42:0],in12[63:43]}) & {in18[20:0],in18[63:21]});
    assign out[1471:1408] = {in12[42:0],in12[63:43]} ^ (~({in18[20:0],in18[63:21]}) & {in24[13:0],in24[63:14]});
    assign out[1407:1344] = {in18[20:0],in18[63:21]} ^ (~({in24[13:0],in24[63:14]}) & in0);
    assign out[1343:1280] = {in24[13:0],in24[63:14]} ^ (~(in0)                      & {in6 [43:0],in6 [63:44]});
    
    assign out[1279:1216] = {in3 [27:0],in3 [63:28]} ^ (~({in9 [19:0],in9 [63:20]}) & {in10[2 :0],in10[63:3 ]});
    assign out[1215:1152] = {in9 [19:0],in9 [63:20]} ^ (~({in10[2 :0],in10[63:3 ]}) & {in16[44:0],in16[63:45]});
    assign out[1151:1088] = {in10[2 :0],in10[63:3 ]} ^ (~({in16[44:0],in16[63:45]}) & {in22[60:0],in22[63:61]});
    assign out[1087:1024] = {in16[44:0],in16[63:45]} ^ (~({in22[60:0],in22[63:61]}) & {in3 [27:0],in3 [63:28]});
    assign out[1023:960 ] = {in22[60:0],in22[63:61]} ^ (~({in3 [27:0],in3 [63:28]}) & {in9 [19:0],in9 [63:20]});
    
    assign out[959 :896 ] = {in1 [0   ],in1 [63:1 ]} ^ (~({in7 [5 :0],in7 [63:6 ]}) & {in13[24:0],in13[63:25]});
    assign out[895 :832 ] = {in7 [5 :0],in7 [63:6 ]} ^ (~({in13[24:0],in13[63:25]}) & {in19[7 :0],in19[63:8 ]});
    assign out[831 :768 ] = {in13[24:0],in13[63:25]} ^ (~({in19[7 :0],in19[63:8 ]}) & {in20[17:0],in20[63:18]});
    assign out[767 :704 ] = {in19[7 :0],in19[63:8 ]} ^ (~({in20[17:0],in20[63:18]}) & {in1 [0   ],in1 [63:1 ]});
    assign out[703 :640 ] = {in20[17:0],in20[63:18]} ^ (~({in1 [0   ],in1 [63:1 ]}) & {in7 [5 :0],in7 [63:6 ]});
    
    assign out[639 :576 ] = {in4 [26:0],in4 [63:27]} ^ (~({in5 [35:0],in5 [63:36]}) & {in11[9 :0],in11[63:10]});
    assign out[575 :512 ] = {in5 [35:0],in5 [63:36]} ^ (~({in11[9 :0],in11[63:10]}) & {in17[14:0],in17[63:15]});
    assign out[511 :448 ] = {in11[9 :0],in11[63:10]} ^ (~({in17[14:0],in17[63:15]}) & {in23[55:0],in23[63:56]});
    assign out[447 :384 ] = {in17[14:0],in17[63:15]} ^ (~({in23[55:0],in23[63:56]}) & {in4 [26:0],in4 [63:27]});
    assign out[383 :320 ] = {in23[55:0],in23[63:56]} ^ (~({in4 [26:0],in4 [63:27]}) & {in5 [35:0],in5 [63:36]});
    
    assign out[319 :256 ] = {in2 [61:0],in2 [63:62]} ^ (~({in8 [54:0],in8 [63:55]}) & {in14[38:0],in14[63:39]});
    assign out[255 :192 ] = {in8 [54:0],in8 [63:55]} ^ (~({in14[38:0],in14[63:39]}) & {in15[40:0],in15[63:41]});
    assign out[191 :128 ] = {in14[38:0],in14[63:39]} ^ (~({in15[40:0],in15[63:41]}) & {in21[1 :0],in21[63:2 ]});
    assign out[127 :64  ] = {in15[40:0],in15[63:41]} ^ (~({in21[1 :0],in21[63:2 ]}) & {in2 [61:0],in2 [63:62]});
    assign out[63  :0   ] = {in21[1 :0],in21[63:2 ]} ^ (~({in2 [61:0],in2 [63:62]}) & {in8 [54:0],in8 [63:55]});

endmodule
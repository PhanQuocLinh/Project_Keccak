`timescale 1ns/1ps
module tb_keccak2stage_ver2 ();
    parameter t = 2;
    parameter DIN_WIDTH  = 1088;
    parameter DOUT_WIDTH = 256;

    wire [DOUT_WIDTH-1:0] out;
    wire hash_ready;
    // wire [4:0] count;
    // wire [1:0] current_state, next_state;
    reg rst_n, clk, first_block, last_block;
    reg [DIN_WIDTH-1:0] IN;
    // wire [1599:0] in_theta, tp_theta, _in_theta, out_iota, w1;
    // wire [7:0] rc;
    initial begin
    clk = 0;
    first_block = 0;
    last_block = 0;
    #t rst_n = 0; 
    // IN = 1088'h0000000048a8ac248000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001;
    // $display("in1_0 = %h", IN);
    #t rst_n = 1; first_block = 1; 
    // start - start
     
    // #(t);
     
    #(1*t);
    IN = 1088'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    $display("in1_0 = %h", IN);
    #(2*t) first_block = 0;
    IN = 1088'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    $display("in2_0 = %h", IN);
    // #(2*t) 
     

    // start - start
    #(47*2*t);
    first_block = 0;
    last_block = 0;
    IN = 1088'h00000000000000000000888888888000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001;
    $display("in1_1 = %h", IN);
    #(2*t);
    last_block  = 1;
    first_block = 0;
    IN = 1088'h00000000000000000000444444448000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001;
    $display("in2_1 = %h", IN);
    #(4*t) first_block = 0; last_block = 0;

    // none - none
    #(47*2*t - t);
    first_block = 1;
    last_block = 0;
    #(t);
    IN = 1088'h0000000048a8ac248000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001;
    $display("in1_0 = %h", IN);
    #(t);
    first_block = 0;
    last_block = 1;
    #(t);
    IN = $random;
    $display("%h", IN);
    #(3*t) last_block = 0;

    #(70*2*t) $stop;
    end

    always @(clk) begin 
        #t clk <= ~clk;
    end

    keccak_2stage_ver2 #(.DIN_WIDTH(DIN_WIDTH), .DOUT_WIDTH(DOUT_WIDTH)) k_2stage 
    (
        .clk(clk),
        .rst_n(rst_n),
        .first_block(first_block),
        .last_block(last_block),
        .in(IN),
        // .count(count),
        .out(out),
        // .current_state(current_state),
        // .next_state(next_state),
        // .in_theta(in_theta),
        // .tp_theta(tp_theta),
        // ._in_theta(_in_theta),
        // .out_iota(out_iota),
        // .w1(w1),
        // .rc(rc),
        .hash_ready(hash_ready)
    );

endmodule






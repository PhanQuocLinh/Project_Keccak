module convert_input_theta(reg1, reg2, reg3, reg4, reg5, reg6, reg7, reg8, reg9, reg10, reg11, reg12, reg13, reg14, reg15, reg16, reg17, reg18, reg19, reg20, reg21 , reg22, reg23, reg24, reg25, in);
    input  [1599:0] in ;
    // input  sel, clk, reset;
    output [63:0 ] reg1;
    output [63:0 ] reg2;
    output [63:0 ] reg3;
    output [63:0 ] reg4;
    output [63:0 ] reg5;
    output [63:0 ] reg6;
    output [63:0 ] reg7;
    output [63:0 ] reg8;
    output [63:0 ] reg9;
    output [63:0 ] reg10;
    output [63:0 ] reg11;
    output [63:0 ] reg12;
    output [63:0 ] reg13;
    output [63:0 ] reg14;
    output [63:0 ] reg15;
    output [63:0 ] reg16;
    output [63:0 ] reg17;
    output [63:0 ] reg18;
    output [63:0 ] reg19;
    output [63:0 ] reg20;
    output [63:0 ] reg21;
    output [63:0 ] reg22;
    output [63:0 ] reg23;
    output [63:0 ] reg24;
    output [63:0 ] reg25;


    assign reg25 = in[63:0];
    assign reg24 = in[127:64];
    assign reg23 = in[191:128];
    assign reg22 = in[255:192];
    assign reg21 = in[319:256];
    assign reg20 = in[383:320];
    assign reg19 = in[447:384];
    assign reg18 = in[511:448];
    assign reg17 = in[575:512];
    assign reg16 = in[639:576];
    assign reg15 = in[703:640];
    assign reg14 = in[767:704];
    assign reg13 = in[831:768];
    assign reg12 = in[895:832];
    assign reg11 = in[959:896];
    assign reg10 = in[1023:960];
    assign reg9 = in[1087:1024];
    assign reg8 = in[1151:1088];
    assign reg7 = in[1215:1152];
    assign reg6 = in[1279:1216];
    assign reg5 = in[1343:1280];
    assign reg4 = in[1407:1344];
    assign reg3 = in[1471:1408];
    assign reg2 = in[1535:1472];
    assign reg1 = in[1599:1536];
endmodule